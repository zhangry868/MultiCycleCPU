library verilog;
use verilog.vl_types.all;
entity Multiple_Cycles_CPU_vlg_tst is
end Multiple_Cycles_CPU_vlg_tst;
